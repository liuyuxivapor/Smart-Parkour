module BZ_bram
#(
    parameter ADDR_WIDTH=11,
    parameter DATA_WIDTH=12
)
(
    input clk,
    input en,
    input [ADDR_WIDTH-1:0] addr_i,
    output reg [DATA_WIDTH-1:0] data_o
);

(*ramstyle="block"*)reg[DATA_WIDTH-1:0]mem[(2**ADDR_WIDTH-1):0] ;

initial 
begin
   $readmemh("E:/ciciec/arm/Smart-Parkour/Software/keil/buzzer_music.hex", mem);
end       
	
always @(posedge clk)
  if (en)
    data_o<=mem[addr_i];

endmodule